`timescale 1ns / 1ps

/*
* FIVE-STAGED PIPELINE DATAPATH
* Description: Implements the 5 pipeline stages: Instruction Fetch (IF),
*              Instruction Decode (ID), Execute (EX), Memory Access (MEM), and Write-Back
*              (WB). Contains the Program Counter (PC), pipeline registers, register file,
*              ALU and data memory. Connects them according to the control
*              signal it receives.
*/

import Pipe_Buf_Reg_PKG::*; // Pipeline register struct definitions

module Datapath #(
    // PARAMETERS
    parameter PC_W = 9,       // Program Counter width.
    parameter INS_W = 32,     // Instruction width.
    parameter RF_ADDRESS = 5, // Register File address width (for 2^5  = 32 registers).
    parameter DATA_W = 32,    // Main Data Path width.
    parameter DM_ADDRESS = 9, // Data Memory address width.
    parameter ALU_CC_W = 4    // ALU Control Code width (for the specific ALU operation).
) (

    // INPUTS
    input logic
    // OBS: Global inputs
    clk,
    reset,

    //OBS2: Control Signals (most are generated by the Controller)
    RegWrite,                                    // Enables writing to the register file.
    ALUsrc,                                      // Selects the ALUS's second operand.
    MemWrite,                                    // Enables writing to the data memory.
    MemRead,                                     // Enables reading from data memory.
    Branch,                                      // Indicates a conditional branch instruction.
    Jump,                                        // Indicates a JAL instruction.
    JumpR,                                       // Indicates a JALT instruction.
    input logic  [          1:0] MemtoReg,       // Selects the data source for register write-back.
    input  logic [          1:0] ALUOp,          // High-level ALU operation category for ALUController.
    input  logic [ALU_CC_W -1:0] ALU_CC,         // specific 4-bit operation code from the ALUController for the ALU.

    // OUTPUTS
    // OBS1: Outputs to the Controller (from decoded instruction).
    output logic [          6:0] opcode,         // The 7-bit opcode of the instruction in the ID stage.
    output logic [          6:0] Funct7,         // The Funct7 field of the instruction in the EX stage.
    output logic [          2:0] Funct3,         // The Funct3 field of the instruction in the EX stage.

    // OBS2: Outputs for verification and debugging (includes OBS3)
    output logic [          1:0] ALUOp_Current,  // The ALUOp for the instruction currently in the EX stage.
    output logic [   DATA_W-1:0] WB_Data,        // The final data being written back to the register file

    // OBS3: Testbench outputs
    output logic [4:0] reg_num,                  // The destination register number in the WB stage.
    output logic [DATA_W-1:0] reg_data,          // The data being written to the register in the WB stage.
    output logic reg_write_sig,                  // The RegWrite signal as seen in the WB stage.
    output logic wr,                             // The MemWrite signal as seen in the MEM stage.
    output logic reade,                          // The MemRead signal as seen in the MEM stage.
    output logic [DM_ADDRESS-1:0] addr,          // The address sent to data memory in the MEM stage.
    output logic [DATA_W-1:0] wr_data,           // The data sent to data memory in the MEM stage.
    output logic [DATA_W-1:0] rd_data            // The data read from data memory in the MEM stage.
);

  // INTERNAL WIRES AND REGISTERS

  // Wires for PC logic
  logic [PC_W-1:0] PC, PCPlus4, Next_PC;

  // Wires for instruction and register data
  logic [INS_W-1:0] Instr;
  logic [DATA_W-1:0] Reg1, Reg2;
  logic [DATA_W-1:0] ReadData;

  // Wires for ALU and Branching
  logic [DATA_W-1:0] SrcB, ALUResult;
  logic [DATA_W-1:0] ExtImm, BrImm, Old_PC_Four, BrPC;
  logic [DATA_W-1:0] WrmuxSrc;
  logic              PcSel; // The master signal to flush pipeline and select new PC.

  // Wires for forwarding logic
  logic [1:0] FAmuxSel;
  logic [1:0] FBmuxSel;
  logic [DATA_W-1:0] FAmux_Result;
  logic [DATA_W-1:0] FBmux_Result;

  // Wire for stalling
  logic Reg_Stall;


  // PIPELINE REGISTER INSTANTIATION
  if_id_reg A;
  id_ex_reg B;
  ex_mem_reg C;
  mem_wb_reg D;

  // -----------------------------
  // STAGE 1: INSTRUCTION FETCH (IF)
  // -----------------------------
  // This stage fetches the next instruction from memory based on the current PC

  // PC + 4 Adder: Calculates the address of the next sequential instruction
  adder #(9) pcadd (
      PC,
      9'b100,
      PCPlus4
  );

  // Next PC Mux: Selects the next value for the PC
  // If PCSel is zero, choose sequential instruction (PC + 4)
  // If PCSel is one, choose the branch/jump target from the BranchUnit (BrPC)
  mux2 #(9) pcmux (
      PCPlus4,
      BrPC[PC_W-1:0],
      PcSel,
      Next_PC
  );

  // PC Register: Stores the current Program Counter. Updates to Next_PC on
  //              each clock edge unless stalled.
  flopr #(9) pcreg (
      clk,
      reset,
      Next_PC,
      Reg_Stall,
      PC
  );

  // Instruction Memory: Fetches the 32-bit instruction from the address
  //                     specified by the PC.
  instructionmemory instr_mem (
      clk,
      PC,
      Instr
  );

  // -----------------------------
  // REGISTER 1: IF/ID (Register A)
  // -----------------------------
  // Latches the fetched instruction and its PC value.

  always @(posedge clk) begin
    if ((reset) || (PcSel))   // If reset or a branch/jump is taken, flush the register
        begin
      A.Curr_Pc <= 0;
      A.Curr_Instr <= 0;
    end
        else if (!Reg_Stall)  // If not stalled, latches the new values.
        begin
      A.Curr_Pc <= PC;
      A.Curr_Instr <= Instr;
    end
    // If stalled, the register holds its current value, creating a bubble.
  end

  // -----------------------------
  // STAGE 2: INSTRUCTION DECODE & REGISTER FETCH (ID)
  // -----------------------------
  // This stage decodes the instruction, reads source register from the Register Fiel, and generates the immediate value.

  // Hazard Detection Unit: Checks for Load-Use hazards
  // Asserts 'Reg_Stall' if a hazard is detected, stalling the pipeline
  HazardDetection detect (
      A.Curr_Instr[19:15],
      A.Curr_Instr[24:20],
      B.rd,
      B.MemRead,
      Reg_Stall
  );

  // Opcode is wired out to the Controller.
  assign opcode = A.Curr_Instr[6:0];

  // Register File: Reads the values from the source register rs1 and rs2
  // OBS: The write operation happens in the WB stage, but the hardware is
  //      described here as a single unit.
  RegFile rf (
      clk,
      reset,
      D.RegWrite,
      D.rd,
      A.Curr_Instr[19:15],
      A.Curr_Instr[24:20],
      WrmuxSrc,
      Reg1,
      Reg2
  );

  // Debugging signals for the Testbench.
  assign reg_num = D.rd;
  assign reg_data = WrmuxSrc;
  assign reg_write_sig = D.RegWrite;

  // Immediate Generator: Decodes the instruction to produce the correct
  //                      sign-extended immediate value.
  imm_Gen Ext_Imm (
      A.Curr_Instr,
      ExtImm
  );

  // -----------------------------
  // REGISTER 2: ID/EX (Register B)
  // -----------------------------
  // Latches all control signals, register values, and the immediate for the EX stage.

  always @(posedge clk) begin
    if ((reset) || (Reg_Stall) || (PcSel))        // If reset, stall, or branch, flushes the register.
        begin
      B.ALUSrc <= 0;
      B.MemtoReg <= 2'b00;
      B.RegWrite <= 0;
      B.MemRead <= 0;
      B.MemWrite <= 0;
      B.ALUOp <= 0;
      B.Branch <= 0;
      B.Jump <= 0;
      B.JumpR <= 0;
      B.Curr_Pc <= 0;
      B.RD_One <= 0;
      B.RD_Two <= 0;
      B.RS_One <= 0;
      B.RS_Two <= 0;
      B.rd <= 0;
      B.ImmG <= 0;
      B.func3 <= 0;
      B.func7 <= 0;
      B.Curr_Instr <= A.Curr_Instr;  //debug tmp
    end else begin                                // Normal operation: latches values from ID stage.
      B.ALUSrc <= ALUsrc;
      B.MemtoReg <= MemtoReg;
      B.RegWrite <= RegWrite;
      B.MemRead <= MemRead;
      B.MemWrite <= MemWrite;
      B.ALUOp <= ALUOp;
      B.Branch <= Branch;
      B.Jump <= Jump;
      B.JumpR <= JumpR;
      B.Curr_Pc <= A.Curr_Pc;
      B.RD_One <= Reg1;
      B.RD_Two <= Reg2;
      B.RS_One <= A.Curr_Instr[19:15];
      B.RS_Two <= A.Curr_Instr[24:20];
      B.rd <= A.Curr_Instr[11:7];
      B.ImmG <= ExtImm;
      B.func3 <= A.Curr_Instr[14:12];
      B.func7 <= A.Curr_Instr[31:25];
      B.Curr_Instr <= A.Curr_Instr;  //debug tmp
    end
  end

  // -----------------------------
  // STAGE 3: EXECUTE (EX)
  // -----------------------------
  // This stage performs the main calculation using the ALU and determines branch/jump outcomes.

  // Forwarding Unit: Resolves data hazards by forwarding results from later
  //                  stages back to the ALU inputs, avoiding stalls.
  ForwardingUnit forunit (
      B.RS_One,
      B.RS_Two,
      C.rd,
      D.rd,
      C.RegWrite,
      D.RegWrite,
      FAmuxSel,
      FBmuxSel
  );

  // Outputs to the ALUController
  assign Funct7 = B.func7;
  assign Funct3 = B.func3;
  assign ALUOp_Current = B.ALUOp;

  // Forwarding Mux for SrcA: Selects first ALU operand
  // Can be from RegFile, MEM stage (C.Alu_Result), or WB stage (WrmuxSrc)
  mux4 #(32) FAmux (
      B.RD_One,
      WrmuxSrc,
      C.Alu_Result,
      B.RD_One,
      FAmuxSel,
      FAmux_Result
  );

  // Forwarding Mux for SrcB: Selects the second register operand
  mux4 #(32) FBmux (
      B.RD_Two,
      WrmuxSrc,
      C.Alu_Result,
      B.RD_Two,
      FBmuxSel,
      FBmux_Result
  );

  // ALU source Mux for SrcB: Chooses between the register operand (from FBmux) or the immediate value, based on the ALUSrc control signal.
  mux2 #(32) srcbmux (
      FBmux_Result,
      B.ImmG,
      B.ALUSrc,
      SrcB
  );

  // ALU: Performs the arithmetic/logical operation
  alu alu_module (
      FAmux_Result,
      SrcB,
      ALU_CC,
      ALUResult
  );

  // Branch Unit: Calculates branch/jump targets and determines if the PC
  //              should be updated
  BranchUnit #(9) brunit (
      B.Curr_Pc,
      B.ImmG,
      B.Branch,
      B.Jump,
      B.JumpR,
      ALUResult,
      BrImm,
      Old_PC_Four,
      BrPC,
      PcSel
  );

  // -----------------------------
  // REGISTER 3: EX/MEM (Register C)
  // -----------------------------
  // Latches the ALU result, data to be stored, and control signals for the MEM stage

  always @(posedge clk) begin
    if (reset)                  // If reset, flushes the register.
        begin
      C.RegWrite <= 0;
      C.MemtoReg <= 2'b00;
      C.MemRead <= 0;
      C.MemWrite <= 0;
      C.Pc_Imm <= 0;
      C.Pc_Four <= 0;
      C.Imm_Out <= 0;
      C.Alu_Result <= 0;
      C.RD_Two <= 0;
      C.rd <= 0;
      C.func3 <= 0;
      C.func7 <= 0;
    end else begin              // Normal operation: latches values from EX stage
      C.RegWrite <= B.RegWrite;
      C.MemtoReg <= B.MemtoReg;
      C.MemRead <= B.MemRead;
      C.MemWrite <= B.MemWrite;
      C.Pc_Imm <= BrImm;
      C.Pc_Four <= Old_PC_Four;
      C.Imm_Out <= B.ImmG;
      C.Alu_Result <= ALUResult;
      C.RD_Two <= FBmux_Result;
      C.rd <= B.rd;
      C.func3 <= B.func3;
      C.func7 <= B.func7;
      C.Curr_Instr <= B.Curr_Instr;  // debug tmp
    end
  end

  // -----------------------------
  // STAGE 4: MEMORY ACCESS (MEM)
  // -----------------------------
  // This stage performs read/write operations to the data memory for LW/SW instructions.
  // For all other instructions, it passes the ALU result through

  // Data Memory Interface: Handles byte-addressable loads and stores
  datamemory data_mem (
      clk,
      C.MemRead,
      C.MemWrite,
      C.Alu_Result[8:0],
      C.RD_Two,
      C.func3,
      ReadData
  );

  // Wire out debugging signals for the testbench
  assign wr = C.MemWrite;
  assign reade = C.MemRead;
  assign addr = C.Alu_Result[8:0];
  assign wr_data = C.RD_Two;
  assign rd_data = ReadData;

  // -----------------------------
  // REGISTER 4: MEM/WB (Register D)
  // -----------------------------
  // Latches the data read from memory and the ALU result for the WB stage

  always @(posedge clk) begin
    if (reset)                      // If reset, flushes registers
        begin
      D.RegWrite <= 0;
      D.MemtoReg <= 2'b00;
      D.Pc_Imm <= 0;
      D.Pc_Four <= 0;
      D.Imm_Out <= 0;
      D.Alu_Result <= 0;
      D.MemReadData <= 0;
      D.rd <= 0;
    end else begin                  // Normal operation: latches values from MEM stage
      D.RegWrite <= C.RegWrite;
      D.MemtoReg <= C.MemtoReg;
      D.Pc_Imm <= C.Pc_Imm;
      D.Pc_Four <= C.Pc_Four;
      D.Imm_Out <= C.Imm_Out;
      D.Alu_Result <= C.Alu_Result;
      D.MemReadData <= ReadData;
      D.rd <= C.rd;
      D.Curr_Instr <= C.Curr_Instr;  //Debug Tmp
    end
  end

  // -----------------------------
  // STAGE 5: WRITE-BACK (WB)
  // -----------------------------
  // This final stage writes the result back into the Register File.

  // Write-Back Mux: Selects the final data to be written to the register file
  // - 2'b00 = From the ALU (For R-Type, I-Type arithmetic)
  // - 2'b01 = From Data Memory (for LW)
  // - 2'b10 = The PC + 4 value (for JAL and JALR)
  mux4 #(32) resmux (
      D.Alu_Result,
      D.MemReadData,
      D.Pc_Four,
      32'hxxxxxxxx,
      D.MemtoReg,
      WrmuxSrc
  );

  // Final output for verification
  assign WB_Data = WrmuxSrc;

endmodule
